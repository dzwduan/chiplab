`ifndef MYCPU_H

    `define MYCPU_H

    `define BR_BUS_WD       33
    `define FS_TO_DS_BUS_WD 64
    `define DS_TO_ES_BUS_WD 151
    `define ES_TO_MS_BUS_WD 72
    `define MS_TO_WS_BUS_WD 70
    `define WS_TO_RF_BUS_WD 38
    // `define ES_TO_DS_FORWARD_BUS 1
    // `define MS_TO_DS_FORWARD_BUS 1

`endif
