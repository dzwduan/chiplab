`include "mycpu.vh"
`default_nettype none
module id_stage (
    input  wire                         clk,
    input  wire                         reset,
    //allowin
    input  wire                         es_allowin,
    output wire                         ds_allowin,
    //from fsF
    input  wire                         fs_to_ds_valid,
    input  wire [`FS_TO_DS_BUS_WD -1:0] fs_to_ds_bus,
    //to es
    output wire                         ds_to_es_valid,
    output wire [`DS_TO_ES_BUS_WD -1:0] ds_to_es_bus,
    //to fs
    output wire [`BR_BUS_WD       -1:0] br_bus,
    //to rf: for write back
    input  wire [`WS_TO_RF_BUS_WD -1:0] ws_to_rf_bus,
    // RAW hazard
    input  wire [`ES_TO_DS_BUS_WD -1:0] es_to_ds_forward_bus,
    input  wire [`MS_TO_DS_BUS_WD -1:0] ms_to_ds_forward_bus,
    input  wire                         es_to_ds_valid,
    input  wire                         ms_to_ds_valid,
    input  wire                         ws_to_ds_valid
);

  wire                        br_taken;
  wire [                31:0] br_target;
  wire [                11:0] alu_op;
  wire                        load_op;
  wire                        store_op;
  wire                        src1_is_pc;
  wire                        src2_is_imm;
  wire                        src2_is_4;
  wire                        res_from_mem;
  wire [                 1:0] mem_size;
  wire                        dst_is_r1;
  wire                        gr_we;
  wire                        src_reg_is_rd;
  wire                        rj_eq_rd;
  wire                        rj_lt_rd_unsign;
  wire                        rj_lt_rd_sign;
  wire [                 4:0] dest;
  wire [                31:0] rj_value;
  wire [                31:0] rkd_value;
  wire [                31:0] ds_imm;
  wire [                 5:0] op_31_26;
  wire [                 3:0] op_25_22;
  wire [                 1:0] op_21_20;
  wire [                 4:0] op_19_15;
  wire [                 4:0] rd;
  wire [                 4:0] rj;
  wire [                 4:0] rk;
  wire [                11:0] i12;
  wire [                19:0] i20;
  wire [                15:0] i16;
  wire [                25:0] i26;

  wire [                63:0] op_31_26_d;
  wire [                15:0] op_25_22_d;
  wire [                 3:0] op_21_20_d;
  wire [                31:0] op_19_15_d;

  wire [                 3:0] mul_div_op;
  wire                        mul_div_sign;

  wire                        inst_add_w;
  wire                        inst_sub_w;
  wire                        inst_slt;
  wire                        inst_slti;
  wire                        inst_sltu;
  wire                        inst_sltui;
  wire                        inst_nor;
  wire                        inst_and;
  wire                        inst_andi;
  wire                        inst_or;
  wire                        inst_ori;
  wire                        inst_xor;
  wire                        inst_xori;
  wire                        inst_sll_w;
  wire                        inst_slli_w;
  wire                        inst_srl_w;
  wire                        inst_srli_w;
  wire                        inst_sra_w;
  wire                        inst_srai_w;
  wire                        inst_addi_w;

  wire                        inst_ld_b;
  wire                        inst_ld_bu;
  wire                        inst_ld_h;
  wire                        inst_ld_hu;
  wire                        inst_ld_w;
  wire                        inst_st_b;
  wire                        inst_st_h;
  wire                        inst_st_w;

  wire                        inst_jirl;
  wire                        inst_b;
  wire                        inst_bl;
  wire                        inst_beq;
  wire                        inst_bne;
  wire                        inst_blt;
  wire                        inst_bge;
  wire                        inst_bltu;
  wire                        inst_bgeu;

  wire                        inst_lu12i_w;
  wire                        inst_mul_w;
  wire                        inst_mulh_w;
  wire                        inst_mulh_wu;
  wire                        inst_div_w;
  wire                        inst_mod_w;
  wire                        inst_div_wu;
  wire                        inst_mod_wu;
  wire                        inst_pcaddu12i;

  wire                        need_ui5;
  wire                        need_ui12;
  wire                        need_si12;
  wire                        need_si16_pc;
  wire                        need_si20;
  wire                        need_si20_pc;
  wire                        need_si26_pc;




  wire                        mem_b_size;
  wire                        mem_h_size;
  wire                        mem_sign_exted;

  wire [                 4:0] rf_raddr1;
  wire [                31:0] rf_rdata1;
  wire [                 4:0] rf_raddr2;
  wire [                31:0] rf_rdata2;
  wire                        rf_we;
  wire [                 4:0] rf_waddr;
  wire [                31:0] rf_wdata;
  reg  [`FS_TO_DS_BUS_WD-1:0] fs_to_ds_bus_r;
  reg                         ds_valid;
  wire [                31:0] ds_pc;
  wire [                31:0] ds_inst;
  wire                        ds_ready_go;
  wire                        inst_need_rj;
  wire                        inst_need_rkd;
  wire                        ms_forward_enable;
  wire [                 4:0] ms_forward_reg;
  wire [                31:0] ms_forward_data;
  wire                        ms_dep_need_stall;
  wire                        es_dep_need_stall;
  wire                        es_forward_enable;
  wire [                 4:0] es_forward_reg;
  wire [                31:0] es_forward_data;
  wire                        rf1_forward_stall;
  wire                        rf2_forward_stall;
  wire                        rf1_es_need_stall;
  wire                        rf2_es_need_stall;
  wire                        rf1_ms_need_stall;
  wire                        rf2_ms_need_stall;
  wire                        rf1_ws_need_stall;
  wire                        rf2_ws_need_stall;




  assign ds_ready_go = ~(rf1_forward_stall || rf2_forward_stall);
  assign ds_allowin = !ds_valid || es_allowin && ds_ready_go;
  assign ds_to_es_valid = ds_valid && ds_ready_go;

  always @(posedge clk) begin
    if (reset || br_taken) begin
      ds_valid <= 1'b0;
    end else if (ds_allowin) begin
      ds_valid <= fs_to_ds_valid;
    end

    if (fs_to_ds_valid && ds_allowin) begin
      fs_to_ds_bus_r <= fs_to_ds_bus;
    end
  end

  assign {ds_pc, ds_inst} = fs_to_ds_bus_r;


  assign op_31_26 = ds_inst[31:26];
  assign op_25_22 = ds_inst[25:22];
  assign op_21_20 = ds_inst[21:20];
  assign op_19_15 = ds_inst[19:15];

  assign rd = ds_inst[4:0];
  assign rj = ds_inst[9:5];
  assign rk = ds_inst[14:10];

  assign i12 = ds_inst[21:10];
  assign i20 = ds_inst[24:5];
  assign i16 = ds_inst[25:10];
  assign i26 = {ds_inst[9:0], ds_inst[25:10]};

  decoder_6_64 u_dec0 (
      .in (op_31_26),
      .out(op_31_26_d)
  );
  decoder_4_16 u_dec1 (
      .in (op_25_22),
      .out(op_25_22_d)
  );
  decoder_2_4 u_dec2 (
      .in (op_21_20),
      .out(op_21_20_d)
  );
  decoder_5_32 u_dec3 (
      .in (op_19_15),
      .out(op_19_15_d)
  );

  assign inst_add_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h00];
  assign inst_sub_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h02];
  assign inst_slt = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h04];
  assign inst_sltu = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h05];
  assign inst_nor = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h08];
  assign inst_and = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h09];
  assign inst_or = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0a];
  assign inst_xor = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0b];
  assign inst_sll_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0e];
  assign inst_srl_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0f];
  assign inst_sra_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h10];
  assign inst_slli_w = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h01];
  assign inst_srli_w = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h09];
  assign inst_srai_w = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h11];
  assign inst_addi_w = op_31_26_d[6'h00] & op_25_22_d[4'ha];

  assign inst_mul_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h18];
  assign inst_mulh_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h19];
  assign inst_mulh_wu = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h1a];
  assign inst_div_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h2] & op_19_15_d[5'h00];
  assign inst_mod_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h2] & op_19_15_d[5'h01];
  assign inst_div_wu = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h2] & op_19_15_d[5'h02];
  assign inst_mod_wu = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h2] & op_19_15_d[5'h03];

  assign inst_slti = op_31_26_d[6'h00] & op_25_22_d[4'h8];
  assign inst_sltui = op_31_26_d[6'h00] & op_25_22_d[4'h9];
  assign inst_addi_w = op_31_26_d[6'h00] & op_25_22_d[4'ha];
  assign inst_andi = op_31_26_d[6'h00] & op_25_22_d[4'hd];
  assign inst_ori = op_31_26_d[6'h00] & op_25_22_d[4'he];
  assign inst_xori = op_31_26_d[6'h00] & op_25_22_d[4'hf];

  assign inst_ld_b = op_31_26_d[6'h0a] & op_25_22_d[4'h0];
  assign inst_ld_h = op_31_26_d[6'h0a] & op_25_22_d[4'h1];
  assign inst_ld_w = op_31_26_d[6'h0a] & op_25_22_d[4'h2];
  assign inst_st_b = op_31_26_d[6'h0a] & op_25_22_d[4'h4];
  assign inst_st_h = op_31_26_d[6'h0a] & op_25_22_d[4'h5];
  assign inst_st_w = op_31_26_d[6'h0a] & op_25_22_d[4'h6];
  assign inst_ld_bu = op_31_26_d[6'h0a] & op_25_22_d[4'h8];
  assign inst_ld_hu = op_31_26_d[6'h0a] & op_25_22_d[4'h9];

  assign inst_jirl = op_31_26_d[6'h13];
  assign inst_b = op_31_26_d[6'h14];
  assign inst_bl = op_31_26_d[6'h15];
  assign inst_beq = op_31_26_d[6'h16];
  assign inst_bne = op_31_26_d[6'h17];
  assign inst_blt = op_31_26_d[6'h18];
  assign inst_bge = op_31_26_d[6'h19];
  assign inst_bltu = op_31_26_d[6'h1a];
  assign inst_bgeu = op_31_26_d[6'h1b];
  assign inst_lu12i_w = op_31_26_d[6'h05] & ~ds_inst[25];
  assign inst_pcaddu12i = op_31_26_d[6'h07] & ~ds_inst[25];

  assign alu_op[0] =inst_add_w      |
                    inst_addi_w     |
                    inst_ld_b       |
                    inst_ld_h       |
                    inst_ld_w       |
                    inst_st_b       |
                    inst_st_h       |
                    inst_st_w       |
                    inst_ld_bu      |
                    inst_ld_hu      |
                    inst_jirl       |
                    inst_bl         |
                    inst_pcaddu12i;



  assign alu_op[1] = inst_sub_w;
  assign alu_op[2] = inst_slt | inst_slti;
  assign alu_op[3] = inst_sltu | inst_sltui;
  assign alu_op[4] = inst_and | inst_andi;
  assign alu_op[5] = inst_nor;
  assign alu_op[6] = inst_or | inst_ori;
  assign alu_op[7] = inst_xor | inst_xori;
  assign alu_op[8] = inst_sll_w | inst_slli_w;
  assign alu_op[9] = inst_srl_w | inst_srli_w;
  assign alu_op[10] = inst_sra_w | inst_srai_w;
  assign alu_op[11] = inst_lu12i_w;

  assign mul_div_op[0] = inst_mul_w;
  assign mul_div_op[1] = inst_mulh_w | inst_mulh_wu;
  assign mul_div_op[2] = inst_div_w | inst_div_wu;
  assign mul_div_op[3] = inst_mod_w | inst_mod_wu;

  assign mul_div_sign = inst_mul_w | inst_mulh_w | inst_div_w | inst_mod_w;

  assign inst_need_rj  =  inst_add_w      |
                        inst_sub_w      |
                        inst_addi_w     |
                        inst_slt        |
                        inst_sltu       |
                        inst_slti       |
                        inst_sltui      |
                        inst_and        |
                        inst_or         |
                        inst_nor        |
                        inst_xor        |
                        inst_andi       |
                        inst_ori        |
                        inst_xori       |
                        inst_mul_w      |
                        inst_mulh_w     |
                        inst_mulh_wu    |
                        inst_div_w      |
                        inst_div_wu     |
                        inst_mod_w      |
                        inst_mod_wu     |
                        inst_sll_w      |
                        inst_srl_w      |
                        inst_sra_w      |
                        inst_slli_w     |
                        inst_srli_w     |
                        inst_srai_w     |
                        inst_beq        |
                        inst_bne        |
                        inst_blt        |
                        inst_bltu       |
                        inst_bge        |
                        inst_bgeu       |
                        inst_jirl       |
                        inst_ld_b       |
                        inst_ld_bu      |
                        inst_ld_h       |
                        inst_ld_hu      |
                        inst_ld_w       |
                        inst_st_b       |
                        inst_st_h       |
                        inst_st_w;


  assign inst_need_rkd = inst_add_w   |
                       inst_sub_w   |
                       inst_slt     |
                       inst_sltu    |
                       inst_and     |
                       inst_or      |
                       inst_nor     |
                       inst_xor     |
                       inst_mul_w   |
                       inst_mulh_w  |
                       inst_mulh_wu |
                       inst_div_w   |
                       inst_div_wu  |
                       inst_mod_w   |
                       inst_mod_wu  |
                       inst_sll_w   |
                       inst_srl_w   |
                       inst_sra_w   |
                       inst_beq     |
                       inst_bne     |
                       inst_blt     |
                       inst_bltu    |
                       inst_bge     |
                       inst_bgeu    |
                       inst_st_b    |
                       inst_st_h    |
                       inst_st_w    ;


  //TODO: dont care pcaddi
  assign need_ui5 = inst_slli_w | inst_srli_w | inst_srai_w;

  assign need_si12     =  inst_addi_w     |
                        inst_ld_b       |
                        inst_ld_h       |
                        inst_ld_w       |
                        inst_st_b       |
                        inst_st_h       |
                        inst_st_w       |
                        inst_ld_bu      |
                        inst_ld_hu      |
                        inst_slti       |
                        inst_sltui      ;

  assign need_ui12 = inst_andi | inst_ori | inst_xori;

  assign need_si16_pc  =  inst_jirl |
                        inst_beq  |
                        inst_bne  |
                        inst_blt  |
                        inst_bge  |
                        inst_bltu |
                        inst_bgeu;

  assign need_si20 = inst_lu12i_w | inst_pcaddu12i;

  assign need_si26_pc = inst_b | inst_bl;

  assign ds_imm = ({32{need_ui5    }} & {27'b0, rk}               ) |
                  ({32{need_si12   }} & {{20{i12[11]}}, i12}      ) |
                  ({32{need_ui12   }} & {20'b0, i12}              ) |
                  ({32{need_si16_pc}} & {{14{i16[15]}}, i16, 2'b0}) |
                  ({32{need_si20}} & {i20, 12'b0})                  |
                  ({32{need_si26_pc}} & {{ 4{i26[25]}}, i26, 2'b0}) ;


  assign src_reg_is_rd = inst_beq | inst_bne | inst_st_w;

  assign src1_is_pc = inst_jirl | inst_bl | inst_pcaddu12i;

  assign src2_is_imm = inst_slli_w     |
                       inst_srli_w     |
                       inst_srai_w     |
                       inst_addi_w     |
                       inst_slti       |
                       inst_sltui      |
                       inst_andi       |
                       inst_ori        |
                       inst_xori       |
                       inst_pcaddu12i  |
                       inst_lu12i_w    |
                       inst_ld_b       |
                       inst_ld_h       |
                       inst_ld_w       |
                       inst_ld_bu      |
                       inst_ld_hu      |
                       inst_st_b       |
                       inst_st_h       |
                       inst_st_w       ;

  assign load_op = inst_ld_b | inst_ld_h | inst_ld_w | inst_ld_bu | inst_ld_hu;
  assign store_op = inst_st_b | inst_st_h | inst_st_w;
  assign mem_b_size = inst_ld_b | inst_ld_bu | inst_st_b;
  assign mem_h_size = inst_ld_h | inst_ld_hu | inst_st_h;
  assign mem_sign_exted = inst_ld_b | inst_ld_h;

  assign mem_size = {mem_h_size, mem_b_size};

  assign res_from_mem = inst_ld_w;
  assign dst_is_r1 = inst_bl;
  assign gr_we =       ~inst_st_b       &
                       ~inst_st_h       &
                       ~inst_st_w       &
                       ~inst_beq        &
                       ~inst_bne        &
                       ~inst_blt        &
                       ~inst_bge        &
                       ~inst_bltu       &
                       ~inst_bgeu       &
                       ~inst_b          ;

  assign dest = dst_is_r1 ? 5'd1 : rd;

  assign rf_raddr1 = rj;
  assign rf_raddr2 = src_reg_is_rd ? rd : rk;

  assign {rf_we,  //37:37
      rf_waddr,  //36:32
      rf_wdata  //31:0
      } = ws_to_rf_bus;

  regfile u_regfile (
      .clk   (clk),
      .raddr1(rf_raddr1),
      .rdata1(rf_rdata1),
      .raddr2(rf_raddr2),
      .rdata2(rf_rdata2),
      .we    (rf_we),
      .waddr (rf_waddr),
      .wdata (rf_wdata)
  );

  assign rj_eq_rd = (rj_value == rkd_value);
  assign rj_lt_rd_unsign = (rj_value < rkd_value);
  assign rj_lt_rd_sign = (rj_value[31] && ~rkd_value[31]) ? 1'b1 :
                         (~rj_value[31] && rkd_value[31]) ? 1'b0 : rj_lt_rd_unsign;

  assign br_taken = (   inst_beq  &&  rj_eq_rd
                    || inst_bne  && !rj_eq_rd
                    || inst_blt  &&  rj_lt_rd_sign
                    || inst_bge  && !rj_lt_rd_sign
                    || inst_bltu &&  rj_lt_rd_unsign
                    || inst_bgeu && !rj_lt_rd_unsign
                    || inst_jirl
                    || inst_bl
                    || inst_b
                  ) && ds_valid;

  assign src2_is_4 = inst_jirl | inst_bl;

  assign br_target = ({32{inst_beq || inst_bne || inst_bl || inst_b ||
                          inst_blt || inst_bge || inst_bltu || inst_bgeu}} & (ds_pc + ds_imm   )) |
                     ({32{inst_jirl}}                                      & (rj_value + ds_imm)) ;


  assign br_bus = {br_taken, br_target};

  assign ds_to_es_bus = {
    mem_sign_exted,  //160:160
    mem_size,  //159:158
    mul_div_op,  //157:154
    mul_div_sign,  //153:153
    alu_op,  //150:139
    load_op,  //138:138
    src1_is_pc,  //137:137
    src2_is_imm,  //136:136
    src2_is_4,  //135:135
    gr_we,  //134:134
    store_op,  //133:133
    dest,  //132:128
    ds_imm,  //127:96
    rj_value,  //95 :64
    rkd_value,  //63 :32
    ds_pc  //31 :0
  };

  // forward path
  assign {es_dep_need_stall,
        es_forward_enable,
        es_forward_reg   ,
        es_forward_data
       } = es_to_ds_forward_bus;

  assign {ms_dep_need_stall,
        ms_forward_enable,
        ms_forward_reg   ,
        ms_forward_data
       } = ms_to_ds_forward_bus;

  assign rf1_es_need_stall = (es_forward_reg == rf_raddr1) && es_forward_enable && inst_need_rj;
  assign rf2_es_need_stall = (es_forward_reg == rf_raddr2) && es_forward_enable && inst_need_rkd;
  assign rf1_ms_need_stall = (ms_forward_reg == rf_raddr1) && ms_forward_enable && inst_need_rj;
  assign rf2_ms_need_stall = (ms_forward_reg == rf_raddr2) && ms_forward_enable && inst_need_rkd;
  assign rf1_ws_need_stall = (rf_waddr == rf_raddr1) && ws_to_ds_valid && inst_need_rj;
  assign rf2_ws_need_stall = (rf_waddr == rf_raddr2) && ws_to_ds_valid && inst_need_rkd;

  assign {rf1_forward_stall, rj_value}  = rf1_es_need_stall ? {es_dep_need_stall, es_forward_data} :
                                          rf1_ms_need_stall ? {ms_dep_need_stall, ms_forward_data} :
                                          rf1_ws_need_stall ? {1'b0, rf_wdata} :
                                                              {1'b0, rf_rdata1};
  assign {rf2_forward_stall, rkd_value} = rf2_es_need_stall ? {es_dep_need_stall, es_forward_data} :
                                          rf2_ms_need_stall ? {ms_dep_need_stall, ms_forward_data} :
                                          rf2_ws_need_stall ? {1'b0, rf_wdata} :
                                                              {1'b0, rf_rdata2};

endmodule
